`timescale 1ns / 1ps

module instr_mem (
    input  logic [31:0] instr_rAddr,
    output logic [31:0] instr_code
);
    logic [31:0] rom[0:63];

    initial begin
        // //R-Type
        // rom[0] =  32'b0000000_00011_00010_000_00101_0110011;  // add  x5, x2, x3
        // rom[1] =  32'b0100000_00011_00010_000_00110_0110011;  // sub  x6, x2, x3
        // rom[2] =  32'b0000000_00011_00010_010_00111_0110011;  // slt  x7, x2, x3
        // rom[3] =  32'b0000000_00011_00010_011_01000_0110011;  // sltu x8, x2, x3
        // rom[4] =  32'b0000000_00011_00010_100_01001_0110011;  // xor  x9, x2, x3
        // rom[5] =  32'b0000000_00011_00010_110_01010_0110011;  // or   x10, x2, x3
        // rom[6] =  32'b0000000_00011_00010_111_01011_0110011;  // and  x11, x2, x3
        // rom[7] =  32'b0000000_00011_00010_001_01100_0110011;  // sll  x12, x2, x3
        // rom[8] =  32'b0000000_00011_00010_101_01101_0110011;  // srl  x13, x2, x3
        // rom[9] =  32'b0100000_00011_00010_101_01110_0110011;  // sra  x14, x2, x3
        // // S-Type
        // rom[10] = 32'b0000000_00100_00000_000_01111_0100011;  // sb  x15, 8(x0)
        // rom[11] = 32'b0000000_00100_00000_001_10000_0100011;  // sh  x16, 8(x0)
        // rom[12] = 32'b0000000_00100_00000_010_10001_0100011;  // sw  x17, 8(x0)
        // //IL_Type
        // rom[13] = 32'b0000000_01100_00010_010_01111_0000011;  // lw   x15, 12(x2)
        // rom[14] = 32'b0000000_01100_00010_001_10000_0000011;  // lh   x16, 12(x2)
        // rom[15] = 32'b0000000_01100_00010_000_10001_0000011;  // lb   x17, 12(x2)
        // rom[16] = 32'b0000000_01100_00010_100_10010_0000011;  // lbu  x18, 12(x2)
        // rom[17] = 32'b0000000_01100_00010_101_10011_0000011;  // lhu  x19, 12(x2)
        // //I_Type_
        // rom[18] = 32'b0000000_01010_00010_000_10100_0010011;  // addi x20, x2, 10
        // rom[19] = 32'b0000000_01010_00010_010_10101_0010011;  // slti x21, x2, 10
        // rom[20] = 32'b0000000_01010_00010_011_10110_0010011;  // sltiu x22, x2, 10
        // rom[21] = 32'b0000000_01010_00010_100_10111_0010011;  // xori x23, x2, 10
        // rom[22] = 32'b0000000_01010_00010_110_11000_0010011;  // ori  x24, x2, 10
        // rom[23] = 32'b0000000_01010_00010_111_11001_0010011;  // andi x25, x2, 10
        // rom[24] = 32'b0000000_00011_00010_001_11010_0010011;  // slli x26, x2, 3
        // rom[25] = 32'b0000000_00011_00010_101_11011_0010011;  // srli x27, x2, 3
        // rom[26] = 32'b0100000_00011_00010_101_11100_0010011;  // srai x28, x2, 3
        //I_Type_test
        // rom[0] =  32'b0000000_01100_00010_010_00100_0000011;  // lw    x4, 12(x2)
        // rom[0] =  32'b0000000_01100_00010_001_00101_0000011;  // lh    x5, 12(x2)
        // rom[2] =  32'b0000000_01100_00010_000_00110_0000011;  // lb    x6, 12(x2)
        // rom[3] =  32'b0000000_01100_00010_100_00111_0000011;  // lbu   x7, 12(x2)
        // rom[4] =  32'b0000000_01100_00010_101_01000_0000011;  // lhu   x8, 12(x2)
        // rom[5] =  32'b0000000_01010_00010_000_01001_0010011;  // addi  x9, x2, 10
        // rom[6] =  32'b0000000_01010_00010_010_01010_0010011;  // slti  x10, x2, 10
        // rom[7] =  32'b0000000_01010_00010_011_01011_0010011;  // sltiu x11, x2, 10
        // rom[8] =  32'b0000000_01010_00010_100_01100_0010011;  // xori  x12, x2, 10
        // rom[9] =  32'b0000000_01010_00010_110_01101_0010011;  // ori   x13, x2, 10
        // rom[10] = 32'b0000000_01010_00010_111_01110_0010011;  // andi  x14, x2, 10
        // rom[11] = 32'b0000000_00011_00010_001_01111_0010011;  // slli  x15, x2, 3
        // rom[12] = 32'b0000000_00011_00010_101_10000_0010011;  // srli  x16, x2, 3
        // rom[13] = 32'b0100000_00011_00010_101_10001_0010011;  // srai  x17, x2, 3
           
        rom [0] = 32'h004182B3; //32'b0000_0000_0100_0001_1000_0010_1011_0011; // add x5, x3, x4
        rom [1] = 32'h409403B3; //32'b0100_0000_1001_0100_0000_0011_1011_0011; // sub x5, x3, x4
        // B_type
        // 32'b0000000_00010_00010_000_10000_1100011;
        // rom[2] = 32'h00_21_08_63; // BEQ x2,x2, 12
        rom[2] = 32'b00000_00000_00000_01100_01000_1110111;
        rom[3] = 32'b00000_00000_00000_01100_01001_1100111;
        // rom[4] = 32'b000000000010_00010_001_10000_1100011;
        // //0010 0001 0101 1000 0 110 0011
        // //0010 0001 0111 10000 1100011
        // rom[5] = 32'h00811323;
        // rom[6] = 32'b000000000010_00010_101_10000_1100011;
        // rom[7] = 32'h00912323;
        // rom[8] = 32'b000000000010_00010_100_10000_1100011;
        // rom[9] = 32'h006103a3;
        // rom[10] = 32'b000000000010_00010_110_10000_1100011;
        // rom[11] = 32'h00C1_2283;
        // rom[12] = 32'b000000000010_00010_111_10000_1100011;
        // rom[13] = 32'h00C3_0413;
        // rom[14] = 32'h00C3_0A93;
    end

    assign instr_code = rom[instr_rAddr[31:2]];

endmodule
